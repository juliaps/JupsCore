module InstructionMemory(AutoClock, Clock, ProgramCounter, Instruction);
	input 	  AutoClock, Clock;
	input 	  [31:0] ProgramCounter;
	output reg [31:0] Instruction;
	reg 		  [31:0] InstMem [512:0];

	always @ (posedge Clock) begin
		
		//main 
		InstMem[0] = 32'b010110_00000_01100_0000000000000000; //loadi r2 0
		InstMem[1] = 32'b001000_00000_01100_0000000000000001; //store r2 r0 1
		InstMem[2] = 32'b010110_00000_01101_0000000000000000; //loadi r3 0
		InstMem[3] = 32'b001000_00000_01101_0000000000000010; //store r3 r0 2
		InstMem[4] = 32'b010110_00000_01110_0000000011011101; //loadi r4 221
		InstMem[5] = 32'b001000_00000_01110_0000000000000011; //store r4 r0 3
		InstMem[6] = 32'b010110_00000_01111_0000000011110011; //loadi r5 243
		InstMem[7] = 32'b001000_00000_01111_0000000000000100; //store r5 r0 4
		InstMem[8] = 32'b010110_00000_10000_0000000000001111; //loadi r6 15
		InstMem[9] = 32'b001000_00000_10000_0000000000000101; //store r6 r0 5
		InstMem[10] = 32'b010110_00000_10001_0000000000110101; //loadi r7 53
		InstMem[11] = 32'b001000_00000_10001_0000000000000110; //store r7 r0 6
		InstMem[12] = 32'b010110_00000_10010_0000000000000001; //loadi r8 1
		InstMem[13] = 32'b001000_00000_10010_0000000000000111; //store r8 r0 7
		InstMem[14] = 32'b000111_00000_11100_0000000000000011; //load r28 r0 3
		InstMem[15] = 32'b000110_11100_00000_11010_00000000000; //mov r26 r28
		InstMem[16] = 32'b011110_11010_11010_11010_00000000000; //exec_proc
		InstMem[17] = 32'b011100_00000_00000_00000_00000000000; //disablereadproc
		InstMem[18] = 32'b011101_00000_00000_00000_00000000000; //disablewriteproc
		InstMem[19] = 32'b000111_00000_10010_0000000000000111; //load r8 r0 7
		InstMem[20] = 32'b010110_00000_10011_0000000000000001; //loadi r9 1
		InstMem[21] = 32'b010001_10011_10010_0000000000111100; //bneq r8 r9 L1
		InstMem[22] = 32'b010000_00000_00010_0000000000111100; //beq t1 r0 L1
		InstMem[23] = 32'b011011_00000_00000_00000_00000000000; //enablereadproc
		InstMem[24] = 32'b000110_11010_00000_00011_00000000000; //mov t2 r26
		InstMem[25] = 32'b000110_11010_00000_11010_00000000000; //mov r26 r26
		InstMem[26] = 32'b011100_00000_00000_00000_00000000000; //disablereadproc
		InstMem[27] = 32'b001000_00000_00011_0000000000000011; //store t2 r0 3
		InstMem[28] = 32'b011011_00000_00000_00000_00000000000; //enablereadproc
		InstMem[29] = 32'b000110_11001_00000_00100_00000000000; //mov t3 r25
		InstMem[30] = 32'b000110_11001_00000_11001_00000000000; //mov r25 r25
		InstMem[31] = 32'b011100_00000_00000_00000_00000000000; //disablereadproc
		InstMem[32] = 32'b001000_00000_00100_0000000000000001; //store t3 r0 1
		InstMem[33] = 32'b000111_00000_11100_0000000000000101; //load r28 r0 5
		InstMem[34] = 32'b011011_00000_00000_00000_00000000000; //enablereadproc
		InstMem[35] = 32'b001000_11100_00000_0000000000000000; //store r0 r28 0
		InstMem[36] = 32'b001000_11100_01011_0000000000000001; //store r1 r28 1
		InstMem[37] = 32'b001000_11100_01100_0000000000000010; //store r2 r28 2
		InstMem[38] = 32'b001000_11100_01101_0000000000000011; //store r3 r28 3
		InstMem[39] = 32'b001000_11100_01110_0000000000000100; //store r4 r28 4
		InstMem[40] = 32'b001000_11100_01111_0000000000000101; //store r5 r28 5
		InstMem[41] = 32'b001000_11100_10000_0000000000000110; //store r6 r28 6
		InstMem[42] = 32'b001000_11100_10001_0000000000000111; //store r7 r28 7
		InstMem[43] = 32'b001000_11100_10010_0000000000001000; //store r8 r28 8
		InstMem[44] = 32'b001000_11100_10011_0000000000001001; //store r9 r28 9
		InstMem[45] = 32'b001000_11100_10100_0000000000001010; //store r10 r28 10
		InstMem[46] = 32'b001000_11100_10101_0000000000001011; //store r11 r28 11
		InstMem[47] = 32'b001000_11100_10110_0000000000001100; //store r12 r28 12
		InstMem[48] = 32'b001000_11100_10111_0000000000001101; //store r13 r28 13
		InstMem[49] = 32'b001000_11100_11000_0000000000001110; //store r14 r28 14
		InstMem[50] = 32'b001000_11100_00000_0000000000001111; //store r15 r28 15
		InstMem[51] = 32'b001000_11100_00000_0000000000010000; //store r16 r28 16
		InstMem[52] = 32'b001000_11100_00000_0000000000010001; //store r17 r28 17
		InstMem[53] = 32'b001000_11100_00000_0000000000010010; //store r18 r28 18
		InstMem[54] = 32'b001000_11100_00000_0000000000010011; //store r19 r28 19
		InstMem[55] = 32'b001000_11100_00000_0000000000010100; //store r20 r28 20
		InstMem[56] = 32'b001000_11100_00000_0000000000010101; //store r21 r28 21
		InstMem[57] = 32'b001000_11100_00000_0000000000010110; //store r22 r28 22
		InstMem[58] = 32'b001000_11100_00000_0000000000010111; //store r23 r28 23
		InstMem[59] = 32'b001000_11100_00000_0000000000011000; //store r24 r28 24
		InstMem[60] = 32'b001000_11100_11001_0000000000011001; //store r25 r28 25
		InstMem[61] = 32'b001000_11100_11010_0000000000011010; //store r26 r28 26
		InstMem[62] = 32'b001000_11100_11011_0000000000011011; //store r27 r28 27
		InstMem[63] = 32'b001000_11100_11100_0000000000011100; //store r28 r28 28
		InstMem[64] = 32'b001000_11100_11101_0000000000011101; //store r29 r28 29
		InstMem[65] = 32'b001000_11100_11110_0000000000011110; //store r30 r28 30
		InstMem[66] = 32'b001000_11100_11111_0000000000011111; //store r31 r28 31
		InstMem[67] = 32'b011100_00000_00000_00000_00000000000; //disablereadproc
		InstMem[68] = 32'b001110_00000_00000_0000000001100011; //j L2
		//label L1
		InstMem[69] = 32'b011011_00000_00000_00000_00000000000; //enablereadproc
		InstMem[70] = 32'b000110_11010_00000_00110_00000000000; //mov t5 r26
		InstMem[71] = 32'b000110_11010_00000_11010_00000000000; //mov r26 r26
		InstMem[72] = 32'b011100_00000_00000_00000_00000000000; //disablereadproc
		InstMem[73] = 32'b001000_00000_00110_0000000000000100; //store t5 r0 4
		InstMem[74] = 32'b011011_00000_00000_00000_00000000000; //enablereadproc
		InstMem[75] = 32'b000110_11001_00000_00111_00000000000; //mov t6 r25
		InstMem[76] = 32'b000110_11001_00000_11001_00000000000; //mov r25 r25
		InstMem[77] = 32'b011100_00000_00000_00000_00000000000; //disablereadproc
		InstMem[78] = 32'b001000_00000_00111_0000000000000010; //store t6 r0 2
		InstMem[79] = 32'b000111_00000_11100_0000000000000110; //load r28 r0 6
		InstMem[80] = 32'b011011_00000_00000_00000_00000000000; //enablereadproc
		InstMem[81] = 32'b001000_11100_00000_0000000000000000; //store r0 r28 0
		InstMem[82] = 32'b001000_11100_01011_0000000000000001; //store r1 r28 1
		InstMem[83] = 32'b001000_11100_01100_0000000000000010; //store r2 r28 2
		InstMem[84] = 32'b001000_11100_01101_0000000000000011; //store r3 r28 3
		InstMem[85] = 32'b001000_11100_01110_0000000000000100; //store r4 r28 4
		InstMem[86] = 32'b001000_11100_01111_0000000000000101; //store r5 r28 5
		InstMem[87] = 32'b001000_11100_10000_0000000000000110; //store r6 r28 6
		InstMem[88] = 32'b001000_11100_10001_0000000000000111; //store r7 r28 7
		InstMem[89] = 32'b001000_11100_10010_0000000000001000; //store r8 r28 8
		InstMem[90] = 32'b001000_11100_10011_0000000000001001; //store r9 r28 9
		InstMem[91] = 32'b001000_11100_10100_0000000000001010; //store r10 r28 10
		InstMem[92] = 32'b001000_11100_10101_0000000000001011; //store r11 r28 11
		InstMem[93] = 32'b001000_11100_10110_0000000000001100; //store r12 r28 12
		InstMem[94] = 32'b001000_11100_10111_0000000000001101; //store r13 r28 13
		InstMem[95] = 32'b001000_11100_11000_0000000000001110; //store r14 r28 14
		InstMem[96] = 32'b001000_11100_00000_0000000000001111; //store r15 r28 15
		InstMem[97] = 32'b001000_11100_00000_0000000000010000; //store r16 r28 16
		InstMem[98] = 32'b001000_11100_00000_0000000000010001; //store r17 r28 17
		InstMem[99] = 32'b001000_11100_00000_0000000000010010; //store r18 r28 18
		InstMem[100] = 32'b001000_11100_00000_0000000000010011; //store r19 r28 19
		InstMem[101] = 32'b001000_11100_00000_0000000000010100; //store r20 r28 20
		InstMem[102] = 32'b001000_11100_00000_0000000000010101; //store r21 r28 21
		InstMem[103] = 32'b001000_11100_00000_0000000000010110; //store r22 r28 22
		InstMem[104] = 32'b001000_11100_00000_0000000000010111; //store r23 r28 23
		InstMem[105] = 32'b001000_11100_00000_0000000000011000; //store r24 r28 24
		InstMem[106] = 32'b001000_11100_11001_0000000000011001; //store r25 r28 25
		InstMem[107] = 32'b001000_11100_11010_0000000000011010; //store r26 r28 26
		InstMem[108] = 32'b001000_11100_11011_0000000000011011; //store r27 r28 27
		InstMem[109] = 32'b001000_11100_11100_0000000000011100; //store r28 r28 28
		InstMem[110] = 32'b001000_11100_11101_0000000000011101; //store r29 r28 29
		InstMem[111] = 32'b001000_11100_11110_0000000000011110; //store r30 r28 30
		InstMem[112] = 32'b001000_11100_11111_0000000000011111; //store r31 r28 31
		InstMem[113] = 32'b011100_00000_00000_00000_00000000000; //disablereadproc
		//label L2
		InstMem[114] = 32'b000111_00000_10111_0000000000000111; //load r13 r0 7
		InstMem[115] = 32'b010110_00000_01011_0000000000000001; //loadi r1 1
		InstMem[116] = 32'b010001_01011_10111_0000000001101110; //bneq r13 r1 L3
		InstMem[117] = 32'b010000_00000_01001_0000000001101110; //beq t8 r0 L3
		InstMem[118] = 32'b000111_00000_01011_0000000000000010; //load r1 r0 2
		InstMem[119] = 32'b010110_00000_01100_0000000000000000; //loadi r2 0
		InstMem[120] = 32'b010001_01100_01011_0000000001101101; //bneq r1 r2 L4
		InstMem[121] = 32'b010000_00000_01010_0000000001101101; //beq t9 r0 L4
		InstMem[122] = 32'b010110_00000_01101_0000000000000010; //loadi r3 2
		InstMem[123] = 32'b001000_00000_01101_0000000000000111; //store r3 r0 7
		//label L4
		InstMem[124] = 32'b001110_00000_00000_0000000001110100; //j L5
		//label L3
		InstMem[125] = 32'b000111_00000_01101_0000000000000001; //load r3 r0 1
		InstMem[126] = 32'b010110_00000_01110_0000000000000000; //loadi r4 0
		InstMem[127] = 32'b010001_01110_01101_0000000001110100; //bneq r3 r4 L6
		InstMem[128] = 32'b010000_00000_00001_0000000001110100; //beq t0 r0 L6
		InstMem[129] = 32'b010110_00000_01111_0000000000000001; //loadi r5 1
		InstMem[130] = 32'b001000_00000_01111_0000000000000111; //store r5 r0 7
		//label L6
		//label L5
		InstMem[131] = 32'b000111_00000_01111_0000000000000111; //load r5 r0 7
		InstMem[132] = 32'b010110_00000_10000_0000000000000001; //loadi r6 1
		InstMem[133] = 32'b010001_10000_01111_0000000010100000; //bneq r5 r6 L7
		InstMem[134] = 32'b010000_00000_00010_0000000010100000; //beq t1 r0 L7
		InstMem[135] = 32'b000111_00000_10000_0000000000000001; //load r6 r0 1
		InstMem[136] = 32'b010110_00000_10001_0000000000000000; //loadi r7 0
		InstMem[137] = 32'b010001_10001_10000_0000000010011111; //bneq r6 r7 L8
		InstMem[138] = 32'b010000_00000_00011_0000000010011111; //beq t2 r0 L8
		InstMem[139] = 32'b000111_00000_11100_0000000000000101; //load r28 r0 5
		InstMem[140] = 32'b011010_00000_00000_00000_00000000000; //enablewriteproc
		InstMem[141] = 32'b000111_11100_00000_0000000000000000; //load r0 r28 0
		InstMem[142] = 32'b000111_11100_01011_0000000000000001; //load r1 r28 1
		InstMem[143] = 32'b000111_11100_01100_0000000000000010; //load r2 r28 2
		InstMem[144] = 32'b000111_11100_01101_0000000000000011; //load r3 r28 3
		InstMem[145] = 32'b000111_11100_01110_0000000000000100; //load r4 r28 4
		InstMem[146] = 32'b000111_11100_01111_0000000000000101; //load r5 r28 5
		InstMem[147] = 32'b000111_11100_10000_0000000000000110; //load r6 r28 6
		InstMem[148] = 32'b000111_11100_10001_0000000000000111; //load r7 r28 7
		InstMem[149] = 32'b000111_11100_10010_0000000000001000; //load r8 r28 8
		InstMem[150] = 32'b000111_11100_10011_0000000000001001; //load r9 r28 9
		InstMem[151] = 32'b000111_11100_10100_0000000000001010; //load r10 r28 10
		InstMem[152] = 32'b000111_11100_10101_0000000000001011; //load r11 r28 11
		InstMem[153] = 32'b000111_11100_10110_0000000000001100; //load r12 r28 12
		InstMem[154] = 32'b000111_11100_10111_0000000000001101; //load r13 r28 13
		InstMem[155] = 32'b000111_11100_11000_0000000000001110; //load r14 r28 14
		InstMem[156] = 32'b000111_11100_00000_0000000000001111; //load r15 r28 15
		InstMem[157] = 32'b000111_11100_00000_0000000000010000; //load r16 r28 16
		InstMem[158] = 32'b000111_11100_00000_0000000000010001; //load r17 r28 17
		InstMem[159] = 32'b000111_11100_00000_0000000000010010; //load r18 r28 18
		InstMem[160] = 32'b000111_11100_00000_0000000000010011; //load r19 r28 19
		InstMem[161] = 32'b000111_11100_00000_0000000000010100; //load r20 r28 20
		InstMem[162] = 32'b000111_11100_00000_0000000000010101; //load r21 r28 21
		InstMem[163] = 32'b000111_11100_00000_0000000000010110; //load r22 r28 22
		InstMem[164] = 32'b000111_11100_00000_0000000000010111; //load r23 r28 23
		InstMem[165] = 32'b000111_11100_00000_0000000000011000; //load r24 r28 24
		InstMem[166] = 32'b000111_11100_11001_0000000000011001; //load r25 r28 25
		InstMem[167] = 32'b000111_11100_11010_0000000000011010; //load r26 r28 26
		InstMem[168] = 32'b000111_11100_11011_0000000000011011; //load r27 r28 27
		InstMem[169] = 32'b000111_11100_11100_0000000000011100; //load r28 r28 28
		InstMem[170] = 32'b000111_11100_11101_0000000000011101; //load r29 r28 29
		InstMem[171] = 32'b000111_11100_11110_0000000000011110; //load r30 r28 30
		InstMem[172] = 32'b000111_11100_11111_0000000000011111; //load r31 r28 31
		InstMem[173] = 32'b011101_00000_00000_00000_00000000000; //disablewriteproc
		InstMem[174] = 32'b000111_00000_11100_0000000000000011; //load r28 r0 3
		InstMem[175] = 32'b000110_11100_00000_11010_00000000000; //mov r26 r28
		InstMem[176] = 32'b011110_11010_11010_11010_00000000000; //exec_proc
		//label L8
		InstMem[177] = 32'b001110_00000_00000_0000000011000111; //j L9
		//label L7
		InstMem[178] = 32'b000111_00000_10001_0000000000000010; //load r7 r0 2
		InstMem[179] = 32'b010110_00000_10010_0000000000000000; //loadi r8 0
		InstMem[180] = 32'b010001_10010_10001_0000000011000111; //bneq r7 r8 L10
		InstMem[181] = 32'b010000_00000_00110_0000000011000111; //beq t5 r0 L10
		InstMem[182] = 32'b000111_00000_11100_0000000000000110; //load r28 r0 6
		InstMem[183] = 32'b011010_00000_00000_00000_00000000000; //enablewriteproc
		InstMem[184] = 32'b000111_11100_00000_0000000000000000; //load r0 r28 0
		InstMem[185] = 32'b000111_11100_01011_0000000000000001; //load r1 r28 1
		InstMem[186] = 32'b000111_11100_01100_0000000000000010; //load r2 r28 2
		InstMem[187] = 32'b000111_11100_01101_0000000000000011; //load r3 r28 3
		InstMem[188] = 32'b000111_11100_01110_0000000000000100; //load r4 r28 4
		InstMem[189] = 32'b000111_11100_01111_0000000000000101; //load r5 r28 5
		InstMem[190] = 32'b000111_11100_10000_0000000000000110; //load r6 r28 6
		InstMem[191] = 32'b000111_11100_10001_0000000000000111; //load r7 r28 7
		InstMem[192] = 32'b000111_11100_10010_0000000000001000; //load r8 r28 8
		InstMem[193] = 32'b000111_11100_10011_0000000000001001; //load r9 r28 9
		InstMem[194] = 32'b000111_11100_10100_0000000000001010; //load r10 r28 10
		InstMem[195] = 32'b000111_11100_10101_0000000000001011; //load r11 r28 11
		InstMem[196] = 32'b000111_11100_10110_0000000000001100; //load r12 r28 12
		InstMem[197] = 32'b000111_11100_10111_0000000000001101; //load r13 r28 13
		InstMem[198] = 32'b000111_11100_11000_0000000000001110; //load r14 r28 14
		InstMem[199] = 32'b000111_11100_00000_0000000000001111; //load r15 r28 15
		InstMem[200] = 32'b000111_11100_00000_0000000000010000; //load r16 r28 16
		InstMem[201] = 32'b000111_11100_00000_0000000000010001; //load r17 r28 17
		InstMem[202] = 32'b000111_11100_00000_0000000000010010; //load r18 r28 18
		InstMem[203] = 32'b000111_11100_00000_0000000000010011; //load r19 r28 19
		InstMem[204] = 32'b000111_11100_00000_0000000000010100; //load r20 r28 20
		InstMem[205] = 32'b000111_11100_00000_0000000000010101; //load r21 r28 21
		InstMem[206] = 32'b000111_11100_00000_0000000000010110; //load r22 r28 22
		InstMem[207] = 32'b000111_11100_00000_0000000000010111; //load r23 r28 23
		InstMem[208] = 32'b000111_11100_00000_0000000000011000; //load r24 r28 24
		InstMem[209] = 32'b000111_11100_11001_0000000000011001; //load r25 r28 25
		InstMem[210] = 32'b000111_11100_11010_0000000000011010; //load r26 r28 26
		InstMem[211] = 32'b000111_11100_11011_0000000000011011; //load r27 r28 27
		InstMem[212] = 32'b000111_11100_11100_0000000000011100; //load r28 r28 28
		InstMem[213] = 32'b000111_11100_11101_0000000000011101; //load r29 r28 29
		InstMem[214] = 32'b000111_11100_11110_0000000000011110; //load r30 r28 30
		InstMem[215] = 32'b000111_11100_11111_0000000000011111; //load r31 r28 31
		InstMem[216] = 32'b011101_00000_00000_00000_00000000000; //disablewriteproc
		InstMem[217] = 32'b000111_00000_11100_0000000000000100; //load r28 r0 4
		InstMem[218] = 32'b000110_11100_00000_11010_00000000000; //mov r26 r28
		InstMem[219] = 32'b011110_11010_11010_11010_00000000000; //exec_proc
		//label L10
		//label L9
		InstMem[220] = 32'b000001_00000_00000_00000_00000000000; //halt

		//main  fatorial
		InstMem[221] = 32'b010110_00000_01100_0000000000000001; //loadi r2 1
		InstMem[222] = 32'b001000_00000_01100_0000000000110000; //store r2 r0 48
		InstMem[223] = 32'b010110_00000_01101_0000000000000101; //loadi r3 5
		InstMem[224] = 32'b001000_00000_01101_0000000000110001; //store r3 r0 49
		InstMem[225] = 32'b010110_00000_01110_0000000000000001; //loadi r4 1
		InstMem[226] = 32'b001000_00000_01110_0000000000110010; //store r4 r0 50
		//label L1
		InstMem[227] = 32'b000111_00000_01110_0000000000110010; //load r4 r0 50
		InstMem[228] = 32'b000111_00000_01111_0000000000110001; //load r5 r0 49
		InstMem[229] = 32'b010010_01110_01111_00001_00000000000; //slt t0 r4 r5
		InstMem[230] = 32'b010000_00000_00001_0000000000010011; //beq t0 r0 L2
		InstMem[231] = 32'b000111_00000_10000_0000000000110010; //load r6 r0 50
		InstMem[232] = 32'b010110_00000_10001_0000000000000001; //loadi r7 1
		InstMem[233] = 32'b000010_10000_10001_00010_00000000000; //add t1 r6 r7
		InstMem[234] = 32'b001000_00000_00010_0000000000110010; //store t1 r0 50
		InstMem[235] = 32'b000111_00000_10010_0000000000110000; //load r8 r0 48
		InstMem[236] = 32'b000111_00000_10011_0000000000110010; //load r9 r0 50
		InstMem[237] = 32'b000100_10010_10011_00011_00000000000; //mult t2 r8 r9
		InstMem[238] = 32'b001000_00000_00011_0000000000110000; //store t2 r0 48
		InstMem[239] = 32'b001110_00000_00000_0000000000000110; //j L1
		//label L2
		InstMem[240] = 32'b000111_00000_11100_0000000000110000; //load r28 r0 48
		InstMem[241] = 32'b001100_11100_00000_00000_00000000000; //out r28
		InstMem[242] = 32'b011001_00000_00000_00000_00000000000; //halt_proc

		//main exponencial
		InstMem[243] = 32'b010110_00000_01100_0000000000000000; //loadi r2 0
		InstMem[244] = 32'b001000_00000_01100_0000000001011001; //store r2 r0 89
		InstMem[245] = 32'b010110_00000_01101_0000000000000001; //loadi r3 1
		InstMem[246] = 32'b001000_00000_01101_0000000001011000; //store r3 r0 88
		InstMem[247] = 32'b010110_00000_01110_0000000000000010; //loadi r4 2
		InstMem[248] = 32'b001000_00000_01110_0000000001010110; //store r4 r0 86
		InstMem[249] = 32'b010110_00000_01111_0000000000001000; //loadi r5 8
		InstMem[250] = 32'b001000_00000_01111_0000000001010111; //store r5 r0 87
		//label L1
		InstMem[251] = 32'b000111_00000_01111_0000000001011001; //load r5 r0 89
		InstMem[252] = 32'b000111_00000_10000_0000000001010111; //load r6 r0 87
		InstMem[253] = 32'b010010_01111_10000_00001_00000000000; //slt t0 r5 r6
		InstMem[254] = 32'b010000_00000_00001_0000000000010101; //beq t0 r0 L2
		InstMem[255] = 32'b000111_00000_10001_0000000001010110; //load r7 r0 86
		InstMem[256] = 32'b000111_00000_10010_0000000001011000; //load r8 r0 88
		InstMem[257] = 32'b000100_10001_10010_00010_00000000000; //mult t1 r7 r8
		InstMem[258] = 32'b001000_00000_00010_0000000001011000; //store t1 r0 88
		InstMem[259] = 32'b000111_00000_10100_0000000001011001; //load r10 r0 89
		InstMem[260] = 32'b010110_00000_10101_0000000000000001; //loadi r11 1
		InstMem[261] = 32'b000010_10100_10101_00011_00000000000; //add t2 r10 r11
		InstMem[262] = 32'b001000_00000_00011_0000000001011001; //store t2 r0 89
		InstMem[263] = 32'b001110_00000_00000_0000000000001000; //j L1
		//label L2
		InstMem[264] = 32'b000111_00000_11100_0000000001011000; //load r28 r0 88
		InstMem[265] = 32'b001100_11100_00000_00000_00000000000; //out r28
		InstMem[266] = 32'b011001_00000_00000_00000_00000000000; //halt_proc

	end
	
	always @ (posedge AutoClock) begin
		Instruction <= InstMem[ProgramCounter];
	end
endmodule