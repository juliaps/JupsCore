module InstructionMemory(AutoClock, Clock, ProgramCounter, Instruction);
	input 	  AutoClock, Clock;
	input 	  [31:0] ProgramCounter;
	output reg [31:0] Instruction;
	reg 		  [31:0] InstMem [99:0];

	always @ (posedge Clock) begin
	
		//InstMem[0] <= 32'b00101100000011100000000000000000; //in r4
		//InstMem[1] <= 32'b01010001110011110000000000000101; //addi r5 r4 5
		//InstMem[2] <= 32'b00110001111000000000000000000000; //out r5
		
		InstMem[0] <= 32'b00011011111000000000000000000000; //mov r0 r31
		InstMem[1] <= 32'b00111000000000000000000000000010; //j main
		//main 
		InstMem[2] <= 32'b00011100000010110000000000000011; //load r1 r0 3
		InstMem[3] <= 32'b01011000000011000000000000000001; //loadi r2 1
		InstMem[4] <= 32'b00100000000011000000000000000011; //store r2 r0 3
		InstMem[5] <= 32'b00101100000000010000000000000000; //in t0
		InstMem[6] <= 32'b00110000001000000000000000000000; //out t0
		InstMem[7] <= 32'b00011100000011000000000000000001; //load r2 r0 1
		InstMem[8] <= 32'b00100000000000010000000000000001; //store t0 r0 1
		InstMem[9] <= 32'b00011100000011010000000000000010; //load r3 r0 2
		InstMem[10] <= 32'b01011000000011100000000000000001; //loadi r4 1
		InstMem[11] <= 32'b00100000000011100000000000000010; //store r4 r0 2
		//label L1
		InstMem[12] <= 32'b00011100000011100000000000000010; //load r4 r0 2
		InstMem[13] <= 32'b00011100000011110000000000000001; //load r5 r0 1
		InstMem[14] <= 32'b01011101110011110001000000000000; //slet t1 r4 r5
		InstMem[15] <= 32'b01000000000000100000000000011011; //beq t1 r0 L2
		InstMem[16] <= 32'b00011100000100000000000000000011; //load r6 r0 3
		InstMem[17] <= 32'b00011100000100010000000000000010; //load r7 r0 2
		InstMem[18] <= 32'b00010010000100010001100000000000; //mult t2 r6 r7
		InstMem[19] <= 32'b00011100000100100000000000000011; //load r8 r0 3
		InstMem[20] <= 32'b00100000000000110000000000000011; //store t2 r0 3
		InstMem[21] <= 32'b00011100000100110000000000000010; //load r9 r0 2
		InstMem[22] <= 32'b01011000000101000000000000000001; //loadi r10 1
		InstMem[23] <= 32'b00001010011101000010000000000000; //add t3 r9 r10
		InstMem[24] <= 32'b00011100000101000000000000000010; //load r10 r0 2
		InstMem[25] <= 32'b00100000000001000000000000000010; //store t3 r0 2
		InstMem[26] <= 32'b00111000000000000000000000001100; //j L1
		//label L2
		InstMem[27] <= 32'b00011100000101010000000000000011; //load r11 r0 3
		InstMem[28] <= 32'b01010011111111110000000000000001; //addi r31 r31 1
		InstMem[29] <= 32'b00100100000111000000000000000000; //push r28
		InstMem[30] <= 32'b00110010101000000000000000000000; //out r11
		InstMem[31] <= 32'b00000100000000000000000000000000; //halt


		
		//MemInst[0] <= 32'b01011000000010110000000000001111; //loadi r1 15
		//MemInst[1] <= 32'b00011100000011000000000000000000; //lw r2 1
		//MemInst[2] <= 32'b00100001100011010000000000000101; //sw r3 r2 5
		//MemInst[3] <= 32'b00011101100011100000000000000101; //lw r4 r2 5
		//MemInst[4] <= 32'b01010001110011110000000000000101; //addi r5 r4 5
		//MemInst[5] <= 32'b01010101110100000000000000000011; //subi r6 r4 3
		//MemInst[6] <= 32'b00110100000000000000000000000000; //jr r0
		


	end
	
	always @ (posedge AutoClock) begin
		Instruction <= InstMem[ProgramCounter];
	end
endmodule