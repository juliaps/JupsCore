module InstructionMemory(AutoClock, Clock, ProgramCounter, Instruction);
	input 	  AutoClock, Clock;
	input 	  [31:0] ProgramCounter;
	output reg [31:0] Instruction;
	reg 		  [31:0] InstMem [799:0];

	always @ (posedge Clock) begin
	
		//InstMem[0] <= 32'b00101100000011100000000000000000; //in r4
		//InstMem[1] <= 32'b01010001110011110000000000000101; //addi r5 r4 5
		//InstMem[2] <= 32'b00110001111000000000000000000000; //out r5
		
		// SO 
		InstMem[0] <= 32'b00011011111000000000000000000000; //mov r0 r31
		InstMem[1] <= 32'b00111000000000000000000000000010; //j main
		//main 
		InstMem[2] <= 32'b00011100000010110000000000001101; //load r1 r0 13
		InstMem[3] <= 32'b01011000000011000000000000000001; //loadi r2 1
		InstMem[4] <= 32'b00100000000011000000000000001101; //store r2 r0 13
		InstMem[5] <= 32'b00011100000011000000000000001001; //load r2 r0 9
		InstMem[6] <= 32'b01011000000011010000000000000011; //loadi r3 3
		InstMem[7] <= 32'b00100000000011010000000000001001; //store r3 r0 9
		InstMem[8] <= 32'b00011100000011010000000000001010; //load r3 r0 10
		InstMem[9] <= 32'b01011000000011100000000000000000; //loadi r4 0
		InstMem[10] <= 32'b00100000000011100000000000001010; //store r4 r0 10
		InstMem[11] <= 32'b00011100000011100000000000000111; //load r4 r0 7
		InstMem[12] <= 32'b01011000000011110000000000000000; //loadi r5 0
		InstMem[13] <= 32'b00100000000011110000000000000111; //store r5 r0 7
		InstMem[14] <= 32'b01011000000110110000000000000000; //loadi r27 0
		InstMem[15] <= 32'b01010011011000010000000000000100; //addi t0 r27 4
		InstMem[16] <= 32'b01011000000011110000001000110100; //loadi r5 564
		InstMem[17] <= 32'b00100000001011110000000000000000; //store r5 t0 0
		InstMem[18] <= 32'b01011000000110110000000000000001; //loadi r27 1
		InstMem[19] <= 32'b01010011011000100000000000000100; //addi t1 r27 4
		InstMem[20] <= 32'b01011000000100000000001001011100; //loadi r6 604
		InstMem[21] <= 32'b00100000010100000000000000000000; //store r6 t1 0
		InstMem[22] <= 32'b01011000000110110000000000000010; //loadi r27 2
		InstMem[23] <= 32'b01010011011000110000000000000100; //addi t2 r27 4
		InstMem[24] <= 32'b01011000000100010000001010010000; //loadi r7 656
		InstMem[25] <= 32'b00100000011100010000000000000000; //store r7 t2 0
		InstMem[26] <= 32'b01011000000110110000000000000000; //loadi r27 0
		InstMem[27] <= 32'b01010011011001000000000000000001; //addi t3 r27 1
		InstMem[28] <= 32'b01011000000100100000000000000000; //loadi r8 0
		InstMem[29] <= 32'b00100000100100100000000000000000; //store r8 t3 0
		InstMem[30] <= 32'b01011000000110110000000000000001; //loadi r27 1
		InstMem[31] <= 32'b01010011011001010000000000000001; //addi t4 r27 1
		InstMem[32] <= 32'b01011000000100110000000000000000; //loadi r9 0
		InstMem[33] <= 32'b00100000101100110000000000000000; //store r9 t4 0
		InstMem[34] <= 32'b01011000000110110000000000000010; //loadi r27 2
		InstMem[35] <= 32'b01010011011001100000000000000001; //addi t5 r27 1
		InstMem[36] <= 32'b01011000000101000000000000000000; //loadi r10 0
		InstMem[37] <= 32'b00100000110101000000000000000000; //store r10 t5 0
		InstMem[38] <= 32'b00011100000010110000000000001000; //load r1 r0 8
		InstMem[39] <= 32'b01011000000011000000000000000000; //loadi r2 0
		InstMem[40] <= 32'b00100000000011000000000000001000; //store r2 r0 8
		//label L1
		InstMem[41] <= 32'b00011100000011000000000000001010; //load r2 r0 10
		InstMem[42] <= 32'b00011100000011010000000000001001; //load r3 r0 9
		InstMem[43] <= 32'b01001001100011010011100000000000; //slt t6 r2 r3
		InstMem[44] <= 32'b01000000000001110000001000011101; //beq t6 r0 L2
		InstMem[45] <= 32'b01011000000111000000000000110010; //loadi r28 50
		InstMem[46] <= 32'b01010011111111110000000000000001; //addi r31 r31 1
		InstMem[47] <= 32'b00100111111111000000000000000000; //push r28 r31 0
		InstMem[48] <= 32'b00101011111111000000000000000000; //pop r28 r31 0
		InstMem[49] <= 32'b01010111111111110000000000000001; //subi r31 r31 1
		InstMem[50] <= 32'b00110011100000000000000000000000; //out r28
		InstMem[51] <= 32'b00011011010010010000000000000000; //mov t8 r26
		InstMem[52] <= 32'b00011100000011100000000000001011; //load r4 r0 11
		InstMem[53] <= 32'b00100000000010010000000000001011; //store t8 r0 11
		InstMem[54] <= 32'b00011100000011110000000000001011; //load r5 r0 11
		InstMem[55] <= 32'b01011000000100000000000000000001; //loadi r6 1
		InstMem[56] <= 32'b01000100000011110000000001010010; //bneq r5 v6 L3
		InstMem[57] <= 32'b01000000000010100000000001010010; //beq t9 r0 L3
		InstMem[58] <= 32'b00011100000110110000000000001000; //load r27 r0 8
		InstMem[59] <= 32'b01010011011000010000000000000001; //addi t0 r27 1
		InstMem[60] <= 32'b01011000000100000000000000000001; //loadi r6 1
		InstMem[61] <= 32'b00100000001100000000000000000000; //store r6 t0 0
		InstMem[62] <= 32'b00011100000100010000000000001010; //load r7 r0 10
		InstMem[63] <= 32'b01011000000100100000000000000001; //loadi r8 1
		InstMem[64] <= 32'b00001010001100100001000000000000; //add t1 r7 r8
		InstMem[65] <= 32'b00011100000100100000000000001010; //load r8 r0 10
		InstMem[66] <= 32'b00100000000000100000000000001010; //store t1 r0 10
		InstMem[67] <= 32'b00011100000100110000000000001101; //load r9 r0 13
		InstMem[68] <= 32'b01011000000101000000000000000001; //loadi r10 1
		InstMem[69] <= 32'b00100000000101000000000000001101; //store r10 r0 13
		InstMem[70] <= 32'b00011100000101000000000000001000; //load r10 r0 8
		InstMem[71] <= 32'b01011000000010110000001110000101; //loadi r1 901
		InstMem[72] <= 32'b00001010100010110001100000000000; //add t2 r10 r1
		InstMem[73] <= 32'b00011100000010110000000000001110; //load r1 r0 14
		InstMem[74] <= 32'b00100000000000110000000000001110; //store t2 r0 14
		InstMem[75] <= 32'b00011100000111000000000000001110; //load r28 r0 14
		InstMem[76] <= 32'b01010011111111110000000000000001; //addi r31 r31 1
		InstMem[77] <= 32'b00100111111111000000000000000000; //push r28 r31 0
		InstMem[78] <= 32'b00101011111111000000000000000000; //pop r28 r31 0
		InstMem[79] <= 32'b01010111111111110000000000000001; //subi r31 r31 1
		InstMem[80] <= 32'b00110011100000000000000000000000; //out r28
		InstMem[81] <= 32'b00111000000000000000000101101010; //j L4
		//label L3
		InstMem[82] <= 32'b00011100000011000000000000001011; //load r2 r0 11
		InstMem[83] <= 32'b01011000000011010000000000000010; //loadi r3 2
		InstMem[84] <= 32'b01000100000011000000000011011111; //bneq r2 v3 L5
		InstMem[85] <= 32'b01000000000001010000000011011111; //beq t4 r0 L5
		InstMem[86] <= 32'b00101100000001100000000000000000; //in t5
		InstMem[87] <= 32'b00110000110000000000000000000000; //out t5
		InstMem[88] <= 32'b00011100000011010000000000001100; //load r3 r0 12
		InstMem[89] <= 32'b00100000000001100000000000001100; //store t5 r0 12
		InstMem[90] <= 32'b00011100000111000000000000001100; //load r28 r0 12
		InstMem[91] <= 32'b01010011111111110000000000000001; //addi r31 r31 1
		InstMem[92] <= 32'b00100111111111000000000000000000; //push r28 r31 0
		InstMem[93] <= 32'b00101011111110000000000000000000; //pop r14 r31 0
		InstMem[94] <= 32'b01010111111111110000000000000001; //subi r31 r31 1
		InstMem[95] <= 32'b01101100000000000000000000000000; //enablewriteproc
		InstMem[96] <= 32'b00011011000110100000000000000000; //mov r26 r14
		InstMem[97] <= 32'b01111000000000000000000000000000; //disablewriteproc
		InstMem[98] <= 32'b00011100000011100000000000001000; //load r4 r0 8
		InstMem[99] <= 32'b01011000000011110000000000000001; //loadi r5 1
		InstMem[100] <= 32'b01000100000011100000000010001000; //bneq r4 v5 L6
		InstMem[101] <= 32'b01000000000010000000000010001000; //beq t7 r0 L6
		InstMem[102] <= 32'b01011000000111000000000000011001; //loadi r28 25
		InstMem[103] <= 32'b01010011111111110000000000000001; //addi r31 r31 1
		InstMem[104] <= 32'b00100111111111000000000000000000; //push r28 r31 0
		InstMem[105] <= 32'b01110000000000000000000000000000; //enablereadproc
		InstMem[106] <= 32'b00100000000000000000000000011001; //store r0 r0 25
		InstMem[107] <= 32'b00100000000010110000000000011010; //store r1 r0 26
		InstMem[108] <= 32'b00100000000011000000000000011011; //store r2 r0 27
		InstMem[109] <= 32'b00100000000011010000000000011100; //store r3 r0 28
		InstMem[110] <= 32'b00100000000011100000000000011101; //store r4 r0 29
		InstMem[111] <= 32'b00100000000011110000000000011110; //store r5 r0 30
		InstMem[112] <= 32'b00100000000100000000000000011111; //store r6 r0 31
		InstMem[113] <= 32'b00100000000100010000000000100000; //store r7 r0 32
		InstMem[114] <= 32'b00100000000100100000000000100001; //store r8 r0 33
		InstMem[115] <= 32'b00100000000100110000000000100010; //store r9 r0 34
		InstMem[116] <= 32'b00100000000101000000000000100011; //store r10 r0 35
		InstMem[117] <= 32'b00100000000101010000000000100100; //store r11 r0 36
		InstMem[118] <= 32'b00100000000101100000000000100101; //store r12 r0 37
		InstMem[119] <= 32'b00100000000101110000000000100110; //store r13 r0 38
		InstMem[120] <= 32'b00100000000110000000000000100111; //store r14 r0 39
		InstMem[121] <= 32'b00100000000110010000000000101000; //store r15 r0 40
		InstMem[122] <= 32'b00100000000000000000000000101001; //store r16 r0 41
		InstMem[123] <= 32'b00100000000000000000000000101010; //store r17 r0 42
		InstMem[124] <= 32'b00100000000000000000000000101011; //store r18 r0 43
		InstMem[125] <= 32'b00100000000000000000000000101100; //store r19 r0 44
		InstMem[126] <= 32'b00100000000000000000000000101101; //store r20 r0 45
		InstMem[127] <= 32'b00100000000000000000000000101110; //store r21 r0 46
		InstMem[128] <= 32'b00100000000000000000000000101111; //store r22 r0 47
		InstMem[129] <= 32'b00100000000000000000000000110000; //store r23 r0 48
		InstMem[130] <= 32'b00100000000000000000000000110001; //store r24 r0 49
		InstMem[131] <= 32'b00100000000000000000000000110010; //store r25 r0 50
		InstMem[132] <= 32'b00100000000110100000000000110011; //store r26 r0 51
		InstMem[133] <= 32'b00100000000110110000000000110100; //store r27 r0 52
		InstMem[134] <= 32'b00100000000111000000000000110101; //store r28 r0 53
		InstMem[135] <= 32'b00100000000111010000000000110110; //store r29 r0 54
		InstMem[136] <= 32'b00100000000111100000000000110111; //store r30 r0 55
		InstMem[137] <= 32'b00100000000111110000000000111000; //store r31 r0 56
		InstMem[138] <= 32'b01110100000000000000000000000000; //disablereadproc
		InstMem[139] <= 32'b00111000000000000000000011010111; //j L7
		//label L6
		InstMem[140] <= 32'b00011100000011110000000000001000; //load r5 r0 8
		InstMem[141] <= 32'b01011000000100000000000000000010; //loadi r6 2
		InstMem[142] <= 32'b01000100000011110000000010110000; //bneq r5 v6 L8
		InstMem[143] <= 32'b01000000000010100000000010110000; //beq t9 r0 L8
		InstMem[144] <= 32'b01011000000111000000000000111111; //loadi r28 63
		InstMem[145] <= 32'b01010011111111110000000000000001; //addi r31 r31 1
		InstMem[146] <= 32'b00100111111111000000000000000000; //push r28 r31 0
		InstMem[147] <= 32'b01110000000000000000000000000000; //enablereadproc
		InstMem[148] <= 32'b00100000000000000000000000111111; //store r0 r0 63
		InstMem[149] <= 32'b00100000000010110000000001000000; //store r1 r0 64
		InstMem[150] <= 32'b00100000000011000000000001000001; //store r2 r0 65
		InstMem[151] <= 32'b00100000000011010000000001000010; //store r3 r0 66
		InstMem[152] <= 32'b00100000000011100000000001000011; //store r4 r0 67
		InstMem[153] <= 32'b00100000000011110000000001000100; //store r5 r0 68
		InstMem[154] <= 32'b00100000000100000000000001000101; //store r6 r0 69
		InstMem[155] <= 32'b00100000000100010000000001000110; //store r7 r0 70
		InstMem[156] <= 32'b00100000000100100000000001000111; //store r8 r0 71
		InstMem[157] <= 32'b00100000000100110000000001001000; //store r9 r0 72
		InstMem[158] <= 32'b00100000000101000000000001001001; //store r10 r0 73
		InstMem[159] <= 32'b00100000000101010000000001001010; //store r11 r0 74
		InstMem[160] <= 32'b00100000000101100000000001001011; //store r12 r0 75
		InstMem[161] <= 32'b00100000000101110000000001001100; //store r13 r0 76
		InstMem[162] <= 32'b00100000000110000000000001001101; //store r14 r0 77
		InstMem[163] <= 32'b00100000000110010000000001001110; //store r15 r0 78
		InstMem[164] <= 32'b00100000000000000000000001001111; //store r16 r0 79
		InstMem[165] <= 32'b00100000000000000000000001010000; //store r17 r0 80
		InstMem[166] <= 32'b00100000000000000000000001010001; //store r18 r0 81
		InstMem[167] <= 32'b00100000000000000000000001010010; //store r19 r0 82
		InstMem[168] <= 32'b00100000000000000000000001010011; //store r20 r0 83
		InstMem[169] <= 32'b00100000000000000000000001010100; //store r21 r0 84
		InstMem[170] <= 32'b00100000000000000000000001010101; //store r22 r0 85
		InstMem[171] <= 32'b00100000000000000000000001010110; //store r23 r0 86
		InstMem[172] <= 32'b00100000000000000000000001010111; //store r24 r0 87
		InstMem[173] <= 32'b00100000000000000000000001011000; //store r25 r0 88
		InstMem[174] <= 32'b00100000000110100000000001011001; //store r26 r0 89
		InstMem[175] <= 32'b00100000000110110000000001011010; //store r27 r0 90
		InstMem[176] <= 32'b00100000000111000000000001011011; //store r28 r0 91
		InstMem[177] <= 32'b00100000000111010000000001011100; //store r29 r0 92
		InstMem[178] <= 32'b00100000000111100000000001011101; //store r30 r0 93
		InstMem[179] <= 32'b00100000000111110000000001011110; //store r31 r0 94
		InstMem[180] <= 32'b01110100000000000000000000000000; //disablereadproc
		InstMem[181] <= 32'b00111000000000000000000011010111; //j L9
		//label L8
		InstMem[182] <= 32'b00011100000100000000000000001000; //load r6 r0 8
		InstMem[183] <= 32'b01011000000100010000000000000011; //loadi r7 3
		InstMem[184] <= 32'b01000100000100000000000011010111; //bneq r6 v7 L10
		InstMem[185] <= 32'b01000000000000100000000011010111; //beq t1 r0 L10
		InstMem[186] <= 32'b01011000000111000000000001100111; //loadi r28 103
		InstMem[187] <= 32'b01010011111111110000000000000001; //addi r31 r31 1
		InstMem[188] <= 32'b00100111111111000000000000000000; //push r28 r31 0
		InstMem[189] <= 32'b01110000000000000000000000000000; //enablereadproc
		InstMem[190] <= 32'b00100000000000000000000001100111; //store r0 r0 103
		InstMem[191] <= 32'b00100000000010110000000001101000; //store r1 r0 104
		InstMem[192] <= 32'b00100000000011000000000001101001; //store r2 r0 105
		InstMem[193] <= 32'b00100000000011010000000001101010; //store r3 r0 106
		InstMem[194] <= 32'b00100000000011100000000001101011; //store r4 r0 107
		InstMem[195] <= 32'b00100000000011110000000001101100; //store r5 r0 108
		InstMem[196] <= 32'b00100000000100000000000001101101; //store r6 r0 109
		InstMem[197] <= 32'b00100000000100010000000001101110; //store r7 r0 110
		InstMem[198] <= 32'b00100000000100100000000001101111; //store r8 r0 111
		InstMem[199] <= 32'b00100000000100110000000001110000; //store r9 r0 112
		InstMem[200] <= 32'b00100000000101000000000001110001; //store r10 r0 113
		InstMem[201] <= 32'b00100000000101010000000001110010; //store r11 r0 114
		InstMem[202] <= 32'b00100000000101100000000001110011; //store r12 r0 115
		InstMem[203] <= 32'b00100000000101110000000001110100; //store r13 r0 116
		InstMem[204] <= 32'b00100000000110000000000001110101; //store r14 r0 117
		InstMem[205] <= 32'b00100000000110010000000001110110; //store r15 r0 118
		InstMem[206] <= 32'b00100000000000000000000001110111; //store r16 r0 119
		InstMem[207] <= 32'b00100000000000000000000001111000; //store r17 r0 120
		InstMem[208] <= 32'b00100000000000000000000001111001; //store r18 r0 121
		InstMem[209] <= 32'b00100000000000000000000001111010; //store r19 r0 122
		InstMem[210] <= 32'b00100000000000000000000001111011; //store r20 r0 123
		InstMem[211] <= 32'b00100000000000000000000001111100; //store r21 r0 124
		InstMem[212] <= 32'b00100000000000000000000001111101; //store r22 r0 125
		InstMem[213] <= 32'b00100000000000000000000001111110; //store r23 r0 126
		InstMem[214] <= 32'b00100000000000000000000001111111; //store r24 r0 127
		InstMem[215] <= 32'b00100000000000000000000010000000; //store r25 r0 128
		InstMem[216] <= 32'b00100000000110100000000010000001; //store r26 r0 129
		InstMem[217] <= 32'b00100000000110110000000010000010; //store r27 r0 130
		InstMem[218] <= 32'b00100000000111000000000010000011; //store r28 r0 131
		InstMem[219] <= 32'b00100000000111010000000010000100; //store r29 r0 132
		InstMem[220] <= 32'b00100000000111100000000010000101; //store r30 r0 133
		InstMem[221] <= 32'b00100000000111110000000010000110; //store r31 r0 134
		InstMem[222] <= 32'b01110100000000000000000000000000; //disablereadproc
		//label L10
		//label L9
		//label L7
		InstMem[223] <= 32'b00011100000110110000000000001000; //load r27 r0 8
		InstMem[224] <= 32'b01010011011001000000000000000100; //addi t3 r27 4
		InstMem[225] <= 32'b00011011001001010000000000000000; //mov t4 r15
		InstMem[226] <= 32'b00100000100001010000000000000000; //store t4 t3 0
		InstMem[227] <= 32'b00011100000100010000000000001101; //load r7 r0 13
		InstMem[228] <= 32'b01011000000100100000000000000001; //loadi r8 1
		InstMem[229] <= 32'b00100000000100100000000000001101; //store r8 r0 13
		InstMem[230] <= 32'b00111000000000000000000101101010; //j L11
		//label L5
		InstMem[231] <= 32'b00011100000100100000000000001011; //load r8 r0 11
		InstMem[232] <= 32'b01011000000100110000000000000011; //loadi r9 3
		InstMem[233] <= 32'b01000100000100100000000101101010; //bneq r8 v9 L12
		InstMem[234] <= 32'b01000000000001100000000101101010; //beq t5 r0 L12
		InstMem[235] <= 32'b00011011000001110000000000000000; //mov t6 r14
		InstMem[236] <= 32'b00011100000100110000000000001100; //load r9 r0 12
		InstMem[237] <= 32'b00100000000001110000000000001100; //store t6 r0 12
		InstMem[238] <= 32'b00011100000111000000000000001100; //load r28 r0 12
		InstMem[239] <= 32'b01010011111111110000000000000001; //addi r31 r31 1
		InstMem[240] <= 32'b00100111111111000000000000000000; //push r28 r31 0
		InstMem[241] <= 32'b00101011111111000000000000000000; //pop r28 r31 0
		InstMem[242] <= 32'b01010111111111110000000000000001; //subi r31 r31 1
		InstMem[243] <= 32'b00110011100000000000000000000000; //out r28
		InstMem[244] <= 32'b00011100000101000000000000001000; //load r10 r0 8
		InstMem[245] <= 32'b01011000000010110000000000000001; //loadi r1 1
		InstMem[246] <= 32'b01000100000101000000000100010100; //bneq r10 v1 L13
		InstMem[247] <= 32'b01000000000010010000000100010100; //beq t8 r0 L13
		InstMem[248] <= 32'b01011000000111000000000000011001; //loadi r28 25
		InstMem[249] <= 32'b01010011111111110000000000000001; //addi r31 r31 1
		InstMem[250] <= 32'b00100111111111000000000000000000; //push r28 r31 0
		InstMem[251] <= 32'b01110000000000000000000000000000; //enablereadproc
		InstMem[252] <= 32'b00100000000000000000000000011001; //store r0 r0 25
		InstMem[253] <= 32'b00100000000010110000000000011010; //store r1 r0 26
		InstMem[254] <= 32'b00100000000011000000000000011011; //store r2 r0 27
		InstMem[255] <= 32'b00100000000011010000000000011100; //store r3 r0 28
		InstMem[256] <= 32'b00100000000011100000000000011101; //store r4 r0 29
		InstMem[257] <= 32'b00100000000011110000000000011110; //store r5 r0 30
		InstMem[258] <= 32'b00100000000100000000000000011111; //store r6 r0 31
		InstMem[259] <= 32'b00100000000100010000000000100000; //store r7 r0 32
		InstMem[260] <= 32'b00100000000100100000000000100001; //store r8 r0 33
		InstMem[261] <= 32'b00100000000100110000000000100010; //store r9 r0 34
		InstMem[262] <= 32'b00100000000101000000000000100011; //store r10 r0 35
		InstMem[263] <= 32'b00100000000101010000000000100100; //store r11 r0 36
		InstMem[264] <= 32'b00100000000101100000000000100101; //store r12 r0 37
		InstMem[265] <= 32'b00100000000101110000000000100110; //store r13 r0 38
		InstMem[266] <= 32'b00100000000110000000000000100111; //store r14 r0 39
		InstMem[267] <= 32'b00100000000110010000000000101000; //store r15 r0 40
		InstMem[268] <= 32'b00100000000000000000000000101001; //store r16 r0 41
		InstMem[269] <= 32'b00100000000000000000000000101010; //store r17 r0 42
		InstMem[270] <= 32'b00100000000000000000000000101011; //store r18 r0 43
		InstMem[271] <= 32'b00100000000000000000000000101100; //store r19 r0 44
		InstMem[272] <= 32'b00100000000000000000000000101101; //store r20 r0 45
		InstMem[273] <= 32'b00100000000000000000000000101110; //store r21 r0 46
		InstMem[274] <= 32'b00100000000000000000000000101111; //store r22 r0 47
		InstMem[275] <= 32'b00100000000000000000000000110000; //store r23 r0 48
		InstMem[276] <= 32'b00100000000000000000000000110001; //store r24 r0 49
		InstMem[277] <= 32'b00100000000000000000000000110010; //store r25 r0 50
		InstMem[278] <= 32'b00100000000110100000000000110011; //store r26 r0 51
		InstMem[279] <= 32'b00100000000110110000000000110100; //store r27 r0 52
		InstMem[280] <= 32'b00100000000111000000000000110101; //store r28 r0 53
		InstMem[281] <= 32'b00100000000111010000000000110110; //store r29 r0 54
		InstMem[282] <= 32'b00100000000111100000000000110111; //store r30 r0 55
		InstMem[283] <= 32'b00100000000111110000000000111000; //store r31 r0 56
		InstMem[284] <= 32'b01110100000000000000000000000000; //disablereadproc
		InstMem[285] <= 32'b00111000000000000000000101100011; //j L14
		//label L13
		InstMem[286] <= 32'b00011100000010110000000000001000; //load r1 r0 8
		InstMem[287] <= 32'b01011000000011000000000000000010; //loadi r2 2
		InstMem[288] <= 32'b01000100000010110000000100111100; //bneq r1 v2 L15
		InstMem[289] <= 32'b01000000000000010000000100111100; //beq t0 r0 L15
		InstMem[290] <= 32'b01011000000111000000000000111111; //loadi r28 63
		InstMem[291] <= 32'b01010011111111110000000000000001; //addi r31 r31 1
		InstMem[292] <= 32'b00100111111111000000000000000000; //push r28 r31 0
		InstMem[293] <= 32'b01110000000000000000000000000000; //enablereadproc
		InstMem[294] <= 32'b00100000000000000000000000111111; //store r0 r0 63
		InstMem[295] <= 32'b00100000000010110000000001000000; //store r1 r0 64
		InstMem[296] <= 32'b00100000000011000000000001000001; //store r2 r0 65
		InstMem[297] <= 32'b00100000000011010000000001000010; //store r3 r0 66
		InstMem[298] <= 32'b00100000000011100000000001000011; //store r4 r0 67
		InstMem[299] <= 32'b00100000000011110000000001000100; //store r5 r0 68
		InstMem[300] <= 32'b00100000000100000000000001000101; //store r6 r0 69
		InstMem[301] <= 32'b00100000000100010000000001000110; //store r7 r0 70
		InstMem[302] <= 32'b00100000000100100000000001000111; //store r8 r0 71
		InstMem[303] <= 32'b00100000000100110000000001001000; //store r9 r0 72
		InstMem[304] <= 32'b00100000000101000000000001001001; //store r10 r0 73
		InstMem[305] <= 32'b00100000000101010000000001001010; //store r11 r0 74
		InstMem[306] <= 32'b00100000000101100000000001001011; //store r12 r0 75
		InstMem[307] <= 32'b00100000000101110000000001001100; //store r13 r0 76
		InstMem[308] <= 32'b00100000000110000000000001001101; //store r14 r0 77
		InstMem[309] <= 32'b00100000000110010000000001001110; //store r15 r0 78
		InstMem[310] <= 32'b00100000000000000000000001001111; //store r16 r0 79
		InstMem[311] <= 32'b00100000000000000000000001010000; //store r17 r0 80
		InstMem[312] <= 32'b00100000000000000000000001010001; //store r18 r0 81
		InstMem[313] <= 32'b00100000000000000000000001010010; //store r19 r0 82
		InstMem[314] <= 32'b00100000000000000000000001010011; //store r20 r0 83
		InstMem[315] <= 32'b00100000000000000000000001010100; //store r21 r0 84
		InstMem[316] <= 32'b00100000000000000000000001010101; //store r22 r0 85
		InstMem[317] <= 32'b00100000000000000000000001010110; //store r23 r0 86
		InstMem[318] <= 32'b00100000000000000000000001010111; //store r24 r0 87
		InstMem[319] <= 32'b00100000000000000000000001011000; //store r25 r0 88
		InstMem[320] <= 32'b00100000000110100000000001011001; //store r26 r0 89
		InstMem[321] <= 32'b00100000000110110000000001011010; //store r27 r0 90
		InstMem[322] <= 32'b00100000000111000000000001011011; //store r28 r0 91
		InstMem[323] <= 32'b00100000000111010000000001011100; //store r29 r0 92
		InstMem[324] <= 32'b00100000000111100000000001011101; //store r30 r0 93
		InstMem[325] <= 32'b00100000000111110000000001011110; //store r31 r0 94
		InstMem[326] <= 32'b01110100000000000000000000000000; //disablereadproc
		InstMem[327] <= 32'b00111000000000000000000101100011; //j L16
		//label L15
		InstMem[328] <= 32'b00011100000011000000000000001000; //load r2 r0 8
		InstMem[329] <= 32'b01011000000011010000000000000011; //loadi r3 3
		InstMem[330] <= 32'b01000100000011000000000101100011; //bneq r2 v3 L17
		InstMem[331] <= 32'b01000000000000110000000101100011; //beq t2 r0 L17
		InstMem[332] <= 32'b01011000000111000000000001100111; //loadi r28 103
		InstMem[333] <= 32'b01010011111111110000000000000001; //addi r31 r31 1
		InstMem[334] <= 32'b00100111111111000000000000000000; //push r28 r31 0
		InstMem[335] <= 32'b01110000000000000000000000000000; //enablereadproc
		InstMem[336] <= 32'b00100000000000000000000001100111; //store r0 r0 103
		InstMem[337] <= 32'b00100000000010110000000001101000; //store r1 r0 104
		InstMem[338] <= 32'b00100000000011000000000001101001; //store r2 r0 105
		InstMem[339] <= 32'b00100000000011010000000001101010; //store r3 r0 106
		InstMem[340] <= 32'b00100000000011100000000001101011; //store r4 r0 107
		InstMem[341] <= 32'b00100000000011110000000001101100; //store r5 r0 108
		InstMem[342] <= 32'b00100000000100000000000001101101; //store r6 r0 109
		InstMem[343] <= 32'b00100000000100010000000001101110; //store r7 r0 110
		InstMem[344] <= 32'b00100000000100100000000001101111; //store r8 r0 111
		InstMem[345] <= 32'b00100000000100110000000001110000; //store r9 r0 112
		InstMem[346] <= 32'b00100000000101000000000001110001; //store r10 r0 113
		InstMem[347] <= 32'b00100000000101010000000001110010; //store r11 r0 114
		InstMem[348] <= 32'b00100000000101100000000001110011; //store r12 r0 115
		InstMem[349] <= 32'b00100000000101110000000001110100; //store r13 r0 116
		InstMem[350] <= 32'b00100000000110000000000001110101; //store r14 r0 117
		InstMem[351] <= 32'b00100000000110010000000001110110; //store r15 r0 118
		InstMem[352] <= 32'b00100000000000000000000001110111; //store r16 r0 119
		InstMem[353] <= 32'b00100000000000000000000001111000; //store r17 r0 120
		InstMem[354] <= 32'b00100000000000000000000001111001; //store r18 r0 121
		InstMem[355] <= 32'b00100000000000000000000001111010; //store r19 r0 122
		InstMem[356] <= 32'b00100000000000000000000001111011; //store r20 r0 123
		InstMem[357] <= 32'b00100000000000000000000001111100; //store r21 r0 124
		InstMem[358] <= 32'b00100000000000000000000001111101; //store r22 r0 125
		InstMem[359] <= 32'b00100000000000000000000001111110; //store r23 r0 126
		InstMem[360] <= 32'b00100000000000000000000001111111; //store r24 r0 127
		InstMem[361] <= 32'b00100000000000000000000010000000; //store r25 r0 128
		InstMem[362] <= 32'b00100000000110100000000010000001; //store r26 r0 129
		InstMem[363] <= 32'b00100000000110110000000010000010; //store r27 r0 130
		InstMem[364] <= 32'b00100000000111000000000010000011; //store r28 r0 131
		InstMem[365] <= 32'b00100000000111010000000010000100; //store r29 r0 132
		InstMem[366] <= 32'b00100000000111100000000010000101; //store r30 r0 133
		InstMem[367] <= 32'b00100000000111110000000010000110; //store r31 r0 134
		InstMem[368] <= 32'b01110100000000000000000000000000; //disablereadproc
		//label L17
		//label L16
		//label L14
		InstMem[369] <= 32'b00011100000110110000000000001000; //load r27 r0 8
		InstMem[370] <= 32'b01010011011001010000000000000100; //addi t4 r27 4
		InstMem[371] <= 32'b00011011001001100000000000000000; //mov t5 r15
		InstMem[372] <= 32'b00100000101001100000000000000000; //store t5 t4 0
		InstMem[373] <= 32'b00011100000011010000000000001101; //load r3 r0 13
		InstMem[374] <= 32'b01011000000011100000000000000001; //loadi r4 1
		InstMem[375] <= 32'b00100000000011100000000000001101; //store r4 r0 13
		//label L12
		//label L11
		//label L4
		InstMem[376] <= 32'b00011100000011100000000000001101; //load r4 r0 13
		InstMem[377] <= 32'b01011000000011110000000000000001; //loadi r5 1
		InstMem[378] <= 32'b01000100000011100000001000011100; //bneq r4 v5 L18
		InstMem[379] <= 32'b01000000000001110000001000011100; //beq t6 r0 L18
		InstMem[380] <= 32'b00011100000011110000000000001000; //load r5 r0 8
		InstMem[381] <= 32'b01011000000100000000000000000001; //loadi r6 1
		InstMem[382] <= 32'b00001001111100000100000000000000; //add t7 r5 r6
		InstMem[383] <= 32'b00011100000100000000000000001000; //load r6 r0 8
		InstMem[384] <= 32'b00100000000010000000000000001000; //store t7 r0 8
		InstMem[385] <= 32'b00011100000100010000000000001000; //load r7 r0 8
		InstMem[386] <= 32'b00011100000100100000000000001001; //load r8 r0 9
		InstMem[387] <= 32'b01000110010100010000000101111010; //bneq r7 r8 L19
		InstMem[388] <= 32'b01000000000010010000000101111010; //beq t8 r0 L19
		InstMem[389] <= 32'b00011100000100110000000000001000; //load r9 r0 8
		InstMem[390] <= 32'b01011000000101000000000000000000; //loadi r10 0
		InstMem[391] <= 32'b00100000000101000000000000001000; //store r10 r0 8
		//label L19
		//label L20
		InstMem[392] <= 32'b00011100000110110000000000001000; //load r27 r0 8
		InstMem[393] <= 32'b01010011011010100000000000000001; //addi t9 r27 1
		InstMem[394] <= 32'b00011101010000010000000000000000; //load t0 t9 0
		InstMem[395] <= 32'b01011000000101000000000000000001; //loadi r10 1
		InstMem[396] <= 32'b01000100000000010000000110001101; //bneq t0 v10 L21
		InstMem[397] <= 32'b01000000000000100000000110001101; //beq t1 r0 L21
		InstMem[398] <= 32'b00011100000101000000000000001000; //load r10 r0 8
		InstMem[399] <= 32'b01011000000010110000000000000001; //loadi r1 1
		InstMem[400] <= 32'b00001010100010110001100000000000; //add t2 r10 r1
		InstMem[401] <= 32'b00011100000010110000000000001000; //load r1 r0 8
		InstMem[402] <= 32'b00100000000000110000000000001000; //store t2 r0 8
		InstMem[403] <= 32'b00011100000011000000000000001000; //load r2 r0 8
		InstMem[404] <= 32'b00011100000011010000000000001001; //load r3 r0 9
		InstMem[405] <= 32'b01000101101011000000000110001100; //bneq r2 r3 L22
		InstMem[406] <= 32'b01000000000001000000000110001100; //beq t3 r0 L22
		InstMem[407] <= 32'b00011100000011100000000000001000; //load r4 r0 8
		InstMem[408] <= 32'b01011000000011110000000000000000; //loadi r5 0
		InstMem[409] <= 32'b00100000000011110000000000001000; //store r5 r0 8
		//label L22
		InstMem[410] <= 32'b00111000000000000000000101111010; //j L20
		//label L21
		InstMem[411] <= 32'b00011100000011110000000000001000; //load r5 r0 8
		InstMem[412] <= 32'b01011000000100000000000000000001; //loadi r6 1
		InstMem[413] <= 32'b01000100000011110000000110110101; //bneq r5 v6 L23
		InstMem[414] <= 32'b01000000000001010000000110110101; //beq t4 r0 L23
		InstMem[415] <= 32'b01011000000111000000000000011001; //loadi r28 25
		InstMem[416] <= 32'b01010011111111110000000000000001; //addi r31 r31 1
		InstMem[417] <= 32'b00100111111111000000000000000000; //push r28 r31 0
		InstMem[418] <= 32'b01101100000000000000000000000000; //enablewriteproc
		InstMem[419] <= 32'b00011100000000000000000000011001; //load r0 r0 25
		InstMem[420] <= 32'b00011100000010110000000000011010; //load r1 r0 26
		InstMem[421] <= 32'b00011100000011000000000000011011; //load r2 r0 27
		InstMem[422] <= 32'b00011100000011010000000000011100; //load r3 r0 28
		InstMem[423] <= 32'b00011100000011100000000000011101; //load r4 r0 29
		InstMem[424] <= 32'b00011100000011110000000000011110; //load r5 r0 30
		InstMem[425] <= 32'b00011100000100000000000000011111; //load r6 r0 31
		InstMem[426] <= 32'b00011100000100010000000000100000; //load r7 r0 32
		InstMem[427] <= 32'b00011100000100100000000000100001; //load r8 r0 33
		InstMem[428] <= 32'b00011100000100110000000000100010; //load r9 r0 34
		InstMem[429] <= 32'b00011100000101000000000000100011; //load r10 r0 35
		InstMem[430] <= 32'b00011100000101010000000000100100; //load r11 r0 36
		InstMem[431] <= 32'b00011100000101100000000000100101; //load r12 r0 37
		InstMem[432] <= 32'b00011100000101110000000000100110; //load r13 r0 38
		InstMem[433] <= 32'b00011100000110000000000000100111; //load r14 r0 39
		InstMem[434] <= 32'b00011100000110010000000000101000; //load r15 r0 40
		InstMem[435] <= 32'b00011100000000000000000000101001; //load r16 r0 41
		InstMem[436] <= 32'b00011100000000000000000000101010; //load r17 r0 42
		InstMem[437] <= 32'b00011100000000000000000000101011; //load r18 r0 43
		InstMem[438] <= 32'b00011100000000000000000000101100; //load r19 r0 44
		InstMem[439] <= 32'b00011100000000000000000000101101; //load r20 r0 45
		InstMem[440] <= 32'b00011100000000000000000000101110; //load r21 r0 46
		InstMem[441] <= 32'b00011100000000000000000000101111; //load r22 r0 47
		InstMem[442] <= 32'b00011100000000000000000000110000; //load r23 r0 48
		InstMem[443] <= 32'b00011100000000000000000000110001; //load r24 r0 49
		InstMem[444] <= 32'b00011100000000000000000000110010; //load r25 r0 50
		InstMem[445] <= 32'b00011100000110100000000000110011; //load r26 r0 51
		InstMem[446] <= 32'b00011100000110110000000000110100; //load r27 r0 52
		InstMem[447] <= 32'b00011100000111000000000000110101; //load r28 r0 53
		InstMem[448] <= 32'b00011100000111010000000000110110; //load r29 r0 54
		InstMem[449] <= 32'b00011100000111100000000000110111; //load r30 r0 55
		InstMem[450] <= 32'b00011100000111110000000000111000; //load r31 r0 56
		InstMem[451] <= 32'b01111000000000000000000000000000; //disablewriteproc
		InstMem[452] <= 32'b00111000000000000000001000000100; //j L24
		//label L23
		InstMem[453] <= 32'b00011100000100000000000000001000; //load r6 r0 8
		InstMem[454] <= 32'b01011000000100010000000000000010; //loadi r7 2
		InstMem[455] <= 32'b01000100000100000000000111011101; //bneq r6 v7 L25
		InstMem[456] <= 32'b01000000000001110000000111011101; //beq t6 r0 L25
		InstMem[457] <= 32'b01011000000111000000000000111111; //loadi r28 63
		InstMem[458] <= 32'b01010011111111110000000000000001; //addi r31 r31 1
		InstMem[459] <= 32'b00100111111111000000000000000000; //push r28 r31 0
		InstMem[460] <= 32'b01101100000000000000000000000000; //enablewriteproc
		InstMem[461] <= 32'b00011100000000000000000000111111; //load r0 r0 63
		InstMem[462] <= 32'b00011100000010110000000001000000; //load r1 r0 64
		InstMem[463] <= 32'b00011100000011000000000001000001; //load r2 r0 65
		InstMem[464] <= 32'b00011100000011010000000001000010; //load r3 r0 66
		InstMem[465] <= 32'b00011100000011100000000001000011; //load r4 r0 67
		InstMem[466] <= 32'b00011100000011110000000001000100; //load r5 r0 68
		InstMem[467] <= 32'b00011100000100000000000001000101; //load r6 r0 69
		InstMem[468] <= 32'b00011100000100010000000001000110; //load r7 r0 70
		InstMem[469] <= 32'b00011100000100100000000001000111; //load r8 r0 71
		InstMem[470] <= 32'b00011100000100110000000001001000; //load r9 r0 72
		InstMem[471] <= 32'b00011100000101000000000001001001; //load r10 r0 73
		InstMem[472] <= 32'b00011100000101010000000001001010; //load r11 r0 74
		InstMem[473] <= 32'b00011100000101100000000001001011; //load r12 r0 75
		InstMem[474] <= 32'b00011100000101110000000001001100; //load r13 r0 76
		InstMem[475] <= 32'b00011100000110000000000001001101; //load r14 r0 77
		InstMem[476] <= 32'b00011100000110010000000001001110; //load r15 r0 78
		InstMem[477] <= 32'b00011100000000000000000001001111; //load r16 r0 79
		InstMem[478] <= 32'b00011100000000000000000001010000; //load r17 r0 80
		InstMem[479] <= 32'b00011100000000000000000001010001; //load r18 r0 81
		InstMem[480] <= 32'b00011100000000000000000001010010; //load r19 r0 82
		InstMem[481] <= 32'b00011100000000000000000001010011; //load r20 r0 83
		InstMem[482] <= 32'b00011100000000000000000001010100; //load r21 r0 84
		InstMem[483] <= 32'b00011100000000000000000001010101; //load r22 r0 85
		InstMem[484] <= 32'b00011100000000000000000001010110; //load r23 r0 86
		InstMem[485] <= 32'b00011100000000000000000001010111; //load r24 r0 87
		InstMem[486] <= 32'b00011100000000000000000001011000; //load r25 r0 88
		InstMem[487] <= 32'b00011100000110100000000001011001; //load r26 r0 89
		InstMem[488] <= 32'b00011100000110110000000001011010; //load r27 r0 90
		InstMem[489] <= 32'b00011100000111000000000001011011; //load r28 r0 91
		InstMem[490] <= 32'b00011100000111010000000001011100; //load r29 r0 92
		InstMem[491] <= 32'b00011100000111100000000001011101; //load r30 r0 93
		InstMem[492] <= 32'b00011100000111110000000001011110; //load r31 r0 94
		InstMem[493] <= 32'b01111000000000000000000000000000; //disablewriteproc
		InstMem[494] <= 32'b00111000000000000000001000000100; //j L26
		//label L25
		InstMem[495] <= 32'b00011100000100010000000000001000; //load r7 r0 8
		InstMem[496] <= 32'b01011000000100100000000000000011; //loadi r8 3
		InstMem[497] <= 32'b01000100000100010000001000000100; //bneq r7 v8 L27
		InstMem[498] <= 32'b01000000000010010000001000000100; //beq t8 r0 L27
		InstMem[499] <= 32'b01011000000111000000000001100111; //loadi r28 103
		InstMem[500] <= 32'b01010011111111110000000000000001; //addi r31 r31 1
		InstMem[501] <= 32'b00100111111111000000000000000000; //push r28 r31 0
		InstMem[502] <= 32'b01101100000000000000000000000000; //enablewriteproc
		InstMem[503] <= 32'b00011100000000000000000001100111; //load r0 r0 103
		InstMem[504] <= 32'b00011100000010110000000001101000; //load r1 r0 104
		InstMem[505] <= 32'b00011100000011000000000001101001; //load r2 r0 105
		InstMem[506] <= 32'b00011100000011010000000001101010; //load r3 r0 106
		InstMem[507] <= 32'b00011100000011100000000001101011; //load r4 r0 107
		InstMem[508] <= 32'b00011100000011110000000001101100; //load r5 r0 108
		InstMem[509] <= 32'b00011100000100000000000001101101; //load r6 r0 109
		InstMem[510] <= 32'b00011100000100010000000001101110; //load r7 r0 110
		InstMem[511] <= 32'b00011100000100100000000001101111; //load r8 r0 111
		InstMem[512] <= 32'b00011100000100110000000001110000; //load r9 r0 112
		InstMem[513] <= 32'b00011100000101000000000001110001; //load r10 r0 113
		InstMem[514] <= 32'b00011100000101010000000001110010; //load r11 r0 114
		InstMem[515] <= 32'b00011100000101100000000001110011; //load r12 r0 115
		InstMem[516] <= 32'b00011100000101110000000001110100; //load r13 r0 116
		InstMem[517] <= 32'b00011100000110000000000001110101; //load r14 r0 117
		InstMem[518] <= 32'b00011100000110010000000001110110; //load r15 r0 118
		InstMem[519] <= 32'b00011100000000000000000001110111; //load r16 r0 119
		InstMem[520] <= 32'b00011100000000000000000001111000; //load r17 r0 120
		InstMem[521] <= 32'b00011100000000000000000001111001; //load r18 r0 121
		InstMem[522] <= 32'b00011100000000000000000001111010; //load r19 r0 122
		InstMem[523] <= 32'b00011100000000000000000001111011; //load r20 r0 123
		InstMem[524] <= 32'b00011100000000000000000001111100; //load r21 r0 124
		InstMem[525] <= 32'b00011100000000000000000001111101; //load r22 r0 125
		InstMem[526] <= 32'b00011100000000000000000001111110; //load r23 r0 126
		InstMem[527] <= 32'b00011100000000000000000001111111; //load r24 r0 127
		InstMem[528] <= 32'b00011100000000000000000010000000; //load r25 r0 128
		InstMem[529] <= 32'b00011100000110100000000010000001; //load r26 r0 129
		InstMem[530] <= 32'b00011100000110110000000010000010; //load r27 r0 130
		InstMem[531] <= 32'b00011100000111000000000010000011; //load r28 r0 131
		InstMem[532] <= 32'b00011100000111010000000010000100; //load r29 r0 132
		InstMem[533] <= 32'b00011100000111100000000010000101; //load r30 r0 133
		InstMem[534] <= 32'b00011100000111110000000010000110; //load r31 r0 134
		InstMem[535] <= 32'b01111000000000000000000000000000; //disablewriteproc
		//label L27
		//label L26
		//label L24
		InstMem[536] <= 32'b00011100000110110000000000001000; //load r27 r0 8
		InstMem[537] <= 32'b01010011011000010000000000000100; //addi t0 r27 4
		InstMem[538] <= 32'b00011100001000100000000000000000; //load t1 t0 0
		InstMem[539] <= 32'b00011000010111000000000000000000; //mov r28 t1
		InstMem[540] <= 32'b01010011111111110000000000000001; //addi r31 r31 1
		InstMem[541] <= 32'b00100111111111000000000000000000; //push r28 r31 0
		InstMem[542] <= 32'b00101011111110010000000000000000; //pop r15 r31 0
		InstMem[543] <= 32'b01010111111111110000000000000001; //subi r31 r31 1
		InstMem[544] <= 32'b00011100000100100000000000001000; //load r8 r0 8
		InstMem[545] <= 32'b01011000000100110000001010111101; //loadi r9 701
		InstMem[546] <= 32'b00001010010100110010000000000000; //add t3 r8 r9
		InstMem[547] <= 32'b00011100000100110000000000001110; //load r9 r0 14
		InstMem[548] <= 32'b00100000000001000000000000001110; //store t3 r0 14
		InstMem[549] <= 32'b00011100000111000000000000001110; //load r28 r0 14
		InstMem[550] <= 32'b01010011111111110000000000000001; //addi r31 r31 1
		InstMem[551] <= 32'b00100111111111000000000000000000; //push r28 r31 0
		InstMem[552] <= 32'b00101011111111000000000000000000; //pop r28 r31 0
		InstMem[553] <= 32'b01010111111111110000000000000001; //subi r31 r31 1
		InstMem[554] <= 32'b00110011100000000000000000000000; //out r28
		InstMem[555] <= 32'b00011100000101000000000000001101; //load r10 r0 13
		InstMem[556] <= 32'b01011000000010110000000000000000; //loadi r1 0
		InstMem[557] <= 32'b00100000000010110000000000001101; //store r1 r0 13
		InstMem[558] <= 32'b01011000000111100000001000110000; //loadi r30 proximo_pc
		InstMem[559] <= 32'b01101000000000000000000000000000; //setprocpc r15 r30
		InstMem[560] <= 32'b01101100000000000000000000000000; //enablewriteproc
		InstMem[561] <= 32'b01110000000000000000000000000000; //enablereadproc
		//label L18
		InstMem[562] <= 32'b00111000000000000000000000101001; //j L1
		//label L2
		InstMem[563] <= 32'b00000100000000000000000000000000; //halt


		// prog1: Fatorial
		InstMem[564] <= 32'b00011011111000000000000000000000; //mov r0 r31
		InstMem[565] <= 32'b00111000000000000000000000000010; //j main
		//main 
		InstMem[566] <= 32'b01111000000000000000000000000000; //disablewriteproc
		InstMem[567] <= 32'b01100100000110100000000000000000; //syscall 2
		InstMem[568] <= 32'b01011000000110010000001000111010; //loadi r15 proximo_pc
		InstMem[569] <= 32'b01111100000000000000000000000000; //setsopc r15 r30
		InstMem[570] <= 32'b00011011010000010000000000000000; //mov t0 r26
		InstMem[571] <= 32'b00011100000010110000000000111011; //load r1 r0 59
		InstMem[572] <= 32'b00100000000000010000000000111011; //store t0 r0 59
		InstMem[573] <= 32'b00011100000011000000000000111100; //load r2 r0 60
		InstMem[574] <= 32'b01011000000011010000000000000001; //loadi r3 1
		InstMem[575] <= 32'b00100000000011010000000000111100; //store r3 r0 60
		//label L1
		InstMem[576] <= 32'b00011100000011010000000000111100; //load r3 r0 60
		InstMem[577] <= 32'b00011100000011100000000000111011; //load r4 r0 59
		InstMem[578] <= 32'b01011101101011100001000000000000; //slet t1 r3 r4
		InstMem[579] <= 32'b01000000000000100000000000011010; //beq t1 r0 L2
		InstMem[580] <= 32'b00011100000011110000000000111010; //load r5 r0 58
		InstMem[581] <= 32'b00011100000100000000000000111100; //load r6 r0 60
		InstMem[582] <= 32'b00010001111100000001100000000000; //mult t2 r5 r6
		InstMem[583] <= 32'b00011100000100010000000000111010; //load r7 r0 58
		InstMem[584] <= 32'b00100000000000110000000000111010; //store t2 r0 58
		InstMem[585] <= 32'b00011100000100100000000000111100; //load r8 r0 60
		InstMem[586] <= 32'b01011000000100110000000000000001; //loadi r9 1
		InstMem[587] <= 32'b00001010010100110010000000000000; //add t3 r8 r9
		InstMem[588] <= 32'b00011100000100110000000000111100; //load r9 r0 60
		InstMem[589] <= 32'b00100000000001000000000000111100; //store t3 r0 60
		InstMem[590] <= 32'b00111000000000000000000000001011; //j L1
		//label L2
		InstMem[591] <= 32'b00011100000111000000000000111010; //load r28 r0 58
		InstMem[592] <= 32'b01010011111111110000000000000001; //addi r31 r31 1
		InstMem[593] <= 32'b00100111111111000000000000000000; //push r28 r31 0
		InstMem[594] <= 32'b01111000000000000000000000000000; //disablewriteproc
		InstMem[595] <= 32'b00101011111110000000000000000000; //pop r14 r31 0
		InstMem[596] <= 32'b01101100000000000000000000000000; //enablewriteproc
		InstMem[597] <= 32'b01010111111111110000000000000001; //subi r31 r31 1
		InstMem[598] <= 32'b01111000000000000000000000000000; //disablewriteproc
		InstMem[599] <= 32'b01100100000110100000000000000000; //syscall 3
		InstMem[600] <= 32'b01011000000110010000001001011010; //loadi r15 proximo_pc
		InstMem[601] <= 32'b01111100000000000000000000000000; //setsopc r15 r30
		InstMem[602] <= 32'b01100100000110100000000000000000; //syscall 1
		InstMem[603] <= 32'b01111100000000000000000000000000; //setsopc r15 r30


		// prog 2 : Fibonnaci
		InstMem[604] <= 32'b00011011111000000000000000000000; //mov r0 r31
		InstMem[605] <= 32'b00111000000000000000000000000010; //j main
		//main 
		InstMem[606] <= 32'b00011100000010110000000001100000; //load r1 r0 96
		InstMem[607] <= 32'b01011000000011000000000000000001; //loadi r2 1
		InstMem[608] <= 32'b00100000000011000000000001100000; //store r2 r0 96
		InstMem[609] <= 32'b00011100000011000000000001100010; //load r2 r0 98
		InstMem[610] <= 32'b01011000000011010000000000000001; //loadi r3 1
		InstMem[611] <= 32'b00100000000011010000000001100010; //store r3 r0 98
		InstMem[612] <= 32'b00011100000011010000000001100011; //load r3 r0 99
		InstMem[613] <= 32'b01011000000011100000000000000001; //loadi r4 1
		InstMem[614] <= 32'b00100000000011100000000001100011; //store r4 r0 99
		InstMem[615] <= 32'b01111000000000000000000000000000; //disablewriteproc
		InstMem[616] <= 32'b01100100000110100000000000000000; //syscall 2
		InstMem[617] <= 32'b01011000000110010000001001101011; //loadi r15 proximo_pc
		InstMem[618] <= 32'b01111100000000000000000000000000; //setsopc r15 r30
		InstMem[619] <= 32'b00011011010000010000000000000000; //mov t0 r26
		InstMem[620] <= 32'b00011100000011100000000001100001; //load r4 r0 97
		InstMem[621] <= 32'b00100000000000010000000001100001; //store t0 r0 97
		//label L1
		InstMem[622] <= 32'b00011100000011110000000001100000; //load r5 r0 96
		InstMem[623] <= 32'b00011100000100000000000001100001; //load r6 r0 97
		InstMem[624] <= 32'b01001001111100000001000000000000; //slt t1 r5 r6
		InstMem[625] <= 32'b01000000000000100000000000101110; //beq t1 r0 L2
		InstMem[626] <= 32'b00011100000111000000000001100010; //load r28 r0 98
		InstMem[627] <= 32'b01010011111111110000000000000001; //addi r31 r31 1
		InstMem[628] <= 32'b00100111111111000000000000000000; //push r28 r31 0
		InstMem[629] <= 32'b01111000000000000000000000000000; //disablewriteproc
		InstMem[630] <= 32'b00101011111110000000000000000000; //pop r14 r31 0
		InstMem[631] <= 32'b01101100000000000000000000000000; //enablewriteproc
		InstMem[632] <= 32'b01010111111111110000000000000001; //subi r31 r31 1
		InstMem[633] <= 32'b01111000000000000000000000000000; //disablewriteproc
		InstMem[634] <= 32'b01100100000110100000000000000000; //syscall 3
		InstMem[635] <= 32'b01011000000110010000001001111101; //loadi r15 proximo_pc
		InstMem[636] <= 32'b01111100000000000000000000000000; //setsopc r15 r30
		InstMem[637] <= 32'b00011100000100010000000001100100; //load r7 r0 100
		InstMem[638] <= 32'b00011100000100100000000001100010; //load r8 r0 98
		InstMem[639] <= 32'b00100000000100100000000001100100; //store r8 r0 100
		InstMem[640] <= 32'b00011100000100110000000001100010; //load r9 r0 98
		InstMem[641] <= 32'b00011100000101000000000001100011; //load r10 r0 99
		InstMem[642] <= 32'b00001010011101000010000000000000; //add t3 r9 r10
		InstMem[643] <= 32'b00011100000101010000000001100010; //load r11 r0 98
		InstMem[644] <= 32'b00100000000001000000000001100010; //store t3 r0 98
		InstMem[645] <= 32'b00011100000101100000000001100011; //load r12 r0 99
		InstMem[646] <= 32'b00011100000101110000000001100100; //load r13 r0 100
		InstMem[647] <= 32'b00100000000101110000000001100011; //store r13 r0 99
		InstMem[648] <= 32'b00011100000110000000000001100000; //load r14 r0 96
		InstMem[649] <= 32'b01011000000010110000000000000001; //loadi r1 1
		InstMem[650] <= 32'b00001011000010110010100000000000; //add t4 r14 r1
		InstMem[651] <= 32'b00011100000010110000000001100000; //load r1 r0 96
		InstMem[652] <= 32'b00100000000001010000000001100000; //store t4 r0 96
		InstMem[653] <= 32'b00111000000000000000000000010001; //j L1
		//label L2
		InstMem[654] <= 32'b01100100000110100000000000000000; //syscall 1
		InstMem[655] <= 32'b01111100000000000000000000000000; //setsopc r15 r30

		// prog 3 : Pontencia
		InstMem[656] <= 32'b00011011111000000000000000000000; //mov r0 r31
		InstMem[657] <= 32'b00111000000000000000000000000010; //j main
		//main 
		InstMem[658] <= 32'b00011100000010110000000010001011; //load r1 r0 139
		InstMem[659] <= 32'b01011000000011000000000000000000; //loadi r2 0
		InstMem[660] <= 32'b00100000000011000000000010001011; //store r2 r0 139
		InstMem[661] <= 32'b00011100000011000000000010001010; //load r2 r0 138
		InstMem[662] <= 32'b01011000000011010000000000000001; //loadi r3 1
		InstMem[663] <= 32'b00100000000011010000000010001010; //store r3 r0 138
		InstMem[664] <= 32'b01111000000000000000000000000000; //disablewriteproc
		InstMem[665] <= 32'b01100100000110100000000000000000; //syscall 2
		InstMem[666] <= 32'b01011000000110010000001010011100; //loadi r15 proximo_pc
		InstMem[667] <= 32'b01111100000000000000000000000000; //setsopc r15 r30
		InstMem[668] <= 32'b00011011010000010000000000000000; //mov t0 r26
		InstMem[669] <= 32'b00011100000011010000000010001000; //load r3 r0 136
		InstMem[670] <= 32'b00100000000000010000000010001000; //store t0 r0 136
		InstMem[671] <= 32'b01111000000000000000000000000000; //disablewriteproc
		InstMem[672] <= 32'b01100100000110100000000000000000; //syscall 2
		InstMem[673] <= 32'b01011000000110010000001010100011; //loadi r15 proximo_pc
		InstMem[674] <= 32'b01111100000000000000000000000000; //setsopc r15 r30
		InstMem[675] <= 32'b00011011010000100000000000000000; //mov t1 r26
		InstMem[676] <= 32'b00011100000011100000000010001001; //load r4 r0 137
		InstMem[677] <= 32'b00100000000000100000000010001001; //store t1 r0 137
		//label L1
		InstMem[678] <= 32'b00011100000011110000000010001011; //load r5 r0 139
		InstMem[679] <= 32'b00011100000100000000000010001001; //load r6 r0 137
		InstMem[680] <= 32'b01001001111100000001100000000000; //slt t2 r5 r6
		InstMem[681] <= 32'b01000000000000110000000000100011; //beq t2 r0 L2
		InstMem[682] <= 32'b00011100000100010000000010001000; //load r7 r0 136
		InstMem[683] <= 32'b00011100000100100000000010001010; //load r8 r0 138
		InstMem[684] <= 32'b00010010001100100010000000000000; //mult t3 r7 r8
		InstMem[685] <= 32'b00011100000100110000000010001010; //load r9 r0 138
		InstMem[686] <= 32'b00100000000001000000000010001010; //store t3 r0 138
		InstMem[687] <= 32'b00011100000101000000000010001011; //load r10 r0 139
		InstMem[688] <= 32'b01011000000101010000000000000001; //loadi r11 1
		InstMem[689] <= 32'b00001010100101010010100000000000; //add t4 r10 r11
		InstMem[690] <= 32'b00011100000101010000000010001011; //load r11 r0 139
		InstMem[691] <= 32'b00100000000001010000000010001011; //store t4 r0 139
		InstMem[692] <= 32'b00111000000000000000000000010100; //j L1
		//label L2
		InstMem[693] <= 32'b00011100000111000000000010001010; //load r28 r0 138
		InstMem[694] <= 32'b01010011111111110000000000000001; //addi r31 r31 1
		InstMem[695] <= 32'b00100111111111000000000000000000; //push r28 r31 0
		InstMem[696] <= 32'b01111000000000000000000000000000; //disablewriteproc
		InstMem[697] <= 32'b00101011111110000000000000000000; //pop r14 r31 0
		InstMem[698] <= 32'b01101100000000000000000000000000; //enablewriteproc
		InstMem[699] <= 32'b01010111111111110000000000000001; //subi r31 r31 1
		InstMem[700] <= 32'b01111000000000000000000000000000; //disablewriteproc
		InstMem[701] <= 32'b01100100000110100000000000000000; //syscall 3
		InstMem[702] <= 32'b01011000000110010000001011000000; //loadi r15 proximo_pc
		InstMem[703] <= 32'b01111100000000000000000000000000; //setsopc r15 r30
		InstMem[704] <= 32'b01100100000110100000000000000000; //syscall 1
		InstMem[705] <= 32'b01111100000000000000000000000000; //setsopc r15 r30


		
		//MemInst[0] <= 32'b01011000000010110000000000001111; //loadi r1 15
		//MemInst[1] <= 32'b00011100000011000000000000000000; //lw r2 1
		//MemInst[2] <= 32'b00100001100011010000000000000101; //sw r3 r2 5
		//MemInst[3] <= 32'b00011101100011100000000000000101; //lw r4 r2 5
		//MemInst[4] <= 32'b01010001110011110000000000000101; //addi r5 r4 5
		//MemInst[5] <= 32'b01010101110100000000000000000011; //subi r6 r4 3
		//MemInst[6] <= 32'b00110100000000000000000000000000; //jr r0
		


	end
	
	always @ (posedge AutoClock) begin
		Instruction <= InstMem[ProgramCounter];
	end
endmodule