module InstructionMemory(AutoClock, Clock, ProgramCounter, Instruction);
	input 	  AutoClock, Clock;
	input 	  [31:0] ProgramCounter;
	output reg [31:0] Instruction;
	reg 		  [31:0] InstMem [799:0];

	always @ (posedge Clock) begin
	
		//InstMem[0] = 32'b00011011111000000000000000000000; //mov r0 r31
		//InstMem[1] = 32'b00010100000000000000000000000000; //j main
		//main 
		//InstMem[2] = 32'b00101100000000010000000000000000; //in t0
		//InstMem[3] = 32'b00110000000000000000100000000000; //out t0
		//InstMem[4] = 32'b00011000000000000000000001000000; //load r1 r0 2
		//InstMem[5] = 32'b00011100000000000000000001000000; //store t0 r0 2
		InstMem[0] = 32'b00000000000000000000000000000000; //load r2 r0 3
		InstMem[1] = 32'b00000000000000000000000000000001; //load r2 r0 3
		InstMem[2] = 32'b00000000000000000000000000000010; //load r2 r0 3
		InstMem[3] = 32'b00000000000000000000000000000011;//load r2 r0 3
		InstMem[4] = 32'b00000000000000000000000000000100; //load r2 r0 3
		InstMem[5] = 32'b00000000000000000000000000000101 ;//load r2 r0 3
		InstMem[6] = 32'b00011000000000000000000001100000; //load r2 r0 3
		InstMem[7] = 32'b01011000000000000000000000100000; //loadi r3 1
		InstMem[8] = 32'b00011100000000000000000001100000; //store r3 r0 3
		//label L1
		InstMem[9] = 32'b00011000000000000000000001100000; //load r3 r0 3
		InstMem[10] = 32'b00011000000000000000000001000000; //load r4 r0 2
		//slet t1
		InstMem[11] = 32'b01000000000000100000000000000000; //beq t1 r0 L2
		InstMem[12] = 32'b00011000000000000000000000100000; //load r5 r0 1
		InstMem[13] = 32'b00011000000000000000000001100000; //load r6 r0 3
		InstMem[14] = 32'b00000001111100000001100000000000; //mult t2 r5 r6
		InstMem[15] = 32'b00011000000000000000000000100000; //load r7 r0 1
		InstMem[16] = 32'b00011100000000000000000000100000; //store t2 r0 1
		InstMem[17] = 32'b00011000000000000000000001100000; //load r8 r0 3
		InstMem[18] = 32'b01011000000000000000000000100000; //loadi r9 1
		InstMem[19] = 32'b00000010010100110010000000000000; //add t3 r8 r9
		InstMem[20] = 32'b00011000000000000000000001100000; //load r9 r0 3
		InstMem[21] = 32'b00011100000000000000000001100000; //store t3 r0 3
		InstMem[22] = 32'b00010100000000000000000000000000; //j L1
		//label L2
		InstMem[23] = 32'b00011000000000000000000000100000; //load r28 r0 1
		InstMem[24] = 32'b00001011111111110000000000000001; //addi r31 r31 1
		InstMem[25] = 32'b00100111111000000000000000000000; //push r28 r31 0
		InstMem[26] = 32'b00101011111111000000000000000000; //pop r28 r31 0
		InstMem[27] = 32'b01010011111111110000000000000001; //subi r31 r31 1
		InstMem[28] = 32'b00110000000000001110000000000000; //out r28
		InstMem[29] = 32'b00000100000000000000000000000000; //halt
		// 

		


	end
	
	always @ (posedge AutoClock) begin
		Instruction <= InstMem[ProgramCounter];
	end
endmodule